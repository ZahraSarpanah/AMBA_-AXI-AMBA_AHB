-------------------------------------------------------------------------------
--
-- Title       : decoder
-- Design      : Amba1
-- Author      : Zahra
-- Company     : A
--
-------------------------------------------------------------------------------
--
-- File        : decode.vhd
-- Generated   : Tue Jan 17 11:43:19 2017
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {decoder} architecture {behavr}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity decoder is
	Haddr : in std_logic_vector(31 downto 0);
	Hselx : out std_logic ;
end decoder;

architecture behavr of decoder is
begin
	

end behavr;
